package timer_ref_pkg;
    localparam FINAL_VALUE = 16;
endpackage