package states_pkg;
    typedef enum bit [1:0] {IDLE, START, DATA, STOP} state_e;
endpackage