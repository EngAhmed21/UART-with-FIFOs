package uart_rx_shared_pkg;
    import states_pkg::*;
    import sys_ref_pkg::*;

    state_e cs_ref;
    bit [SCNT_BIT-1:0] s_cnt_ref;
endpackage