package ref_pkg;
    import states_pkg::*;
    import param_pkg::*;

    state_e cs_ref;
    bit [SCNT_BIT-1:0] s_cnt_ref;
endpackage