package FIFO_ref_pkg;
    localparam WIDTH = 8;
    localparam DEPTH = 128;
endpackage